module buff_coass(input d,en,output y);
assign y= d & en;
endmodule
