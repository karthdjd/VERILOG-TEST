module and_g_lev(input a,input b,output c);
assign c=a&b;
endmodule

