module buff_gl(input d,en,output y);
buf(y,d,en);
endmodule

